`timescale 1ns/1ps

module tb_controller;

	reg clock;
	reg reset;
	reg bist_start;
	reg bist_end_reached;

	wire bist_end;
	wire mode;
	wire init;
	wire running;
	wire finish;

	reg s, dv, l_in;
	reg [1:0] test_in;

	wire cut_fz_L;
	wire cut_lclk;
	wire [4:0] cut_read_a;
	wire [1:0] cut_test_out;
	wire pass_nfail;

	top_module top_inst (
		.clock(clock),
		.reset(reset),
		.bist_start(bist_start),
		.s(s),
		.dv(dv),
		.l_in(l_in),
		.test_in(test_in),
		.pass_nfail(pass_nfail),
		.bist_end(bist_end),
		.cut_fz_L(cut_fz_L),
		.cut_lclk(cut_lclk),
		.cut_read_a(cut_read_a),
		.cut_test_out(cut_test_out)
	);

	always #2000 clock = ~clock;

	always @(posedge clock) begin
		if (bist_end) begin
			$display("t=%0t | reset=%b bist_start=%b | bist_end=%b",
				$time, reset, bist_start, bist_end);
		end
	end

	initial begin
		clock = 1'b0;
		reset = 1'b1;
		bist_start = 1'b0;
		s = 1'b0;
		dv = 1'b0;
		l_in = 1'b0;
		test_in = 2'b00;
		bist_end_reached = 1'b0;

		// Sequence one
		#8000 reset = 0;
		#4000 bist_start = 1;

		begin: loop_block_1
			repeat (20000) begin
				@(posedge clock);
				
				if (bist_end === 1'b1) begin
					$display("=== Controller reached bist_end (Sequence one) ===");
					bist_end_reached = 1;
					disable loop_block_1;
				end
			end
		end

		if (!bist_end_reached) begin
			$display("=== Controller did not reach bist_end (Sequence one) ===");
			$finish;
		end
		#4000 bist_end_reached = 0;

		// Sequence two
		#100 bist_start = 0;
		#4000 bist_start = 1;
		#8000 bist_start = 0;
		#8000 bist_start = 1;
		#4000 reset = 1;
		
		#4000 bist_start = 0;
		#4000 bist_start = 1;
		#4000 reset = 0;
		#4000 bist_start = 0;
		#4000 bist_start = 1;

		begin: loop_block_2
			repeat (20000) begin
				@(posedge clock);
				
				if (bist_end === 1'b1) begin
					$display("=== Controller reached bist_end (Sequence two) ===");
					bist_end_reached = 1;
					disable loop_block_2;
				end
			end
		end

		if (!bist_end_reached) begin
			$display("=== Controller did not reach bist_end (Sequence two) ===");
			$finish;
		end
		#4000 bist_end_reached = 0;

		$finish;
	end
endmodule
